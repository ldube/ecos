# ====================================================================
#
#      hal_mn10300_am33.cdl
#
#      MN10300/AM33 variant architectural HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  nickg
# Contributors:   dmoseley
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MN10300_AM33 {
    display "MN10300 AM33 variant"
    parent        CYGPKG_HAL_MN10300
    implements CYGINT_HAL_MN10300_VARIANT
    hardware
    include_dir   cyg/hal
    define_header hal_mn10300_am33.h
    description   "
           The MN10300 AM33 variant HAL package provides generic
           support for this processor architecture. It is also
           necessary to select a specific target platform HAL
           package."

    cdl_option CYGHWR_HAL_MN10300_AM33_REVISION {
        display       "AM33 architecture revision"
        flavor        data
        calculated {1}
        description   "
            The AM33 architecture revision."
    }

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_mn10300.h>"
    }

    compile       var_misc.c variant.S

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/mn10300_am33.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/mn10300_am33.ld" }
    }

    cdl_option CYGSEM_HAL_UNCACHED_FLASH_ACCESS {
        display       "Caching needn't be disabled to access flash"
        flavor        bool
        default_value 0
        description   "
            Enable this option if the hardware is able to program the flash
            without turning off CPU data caching."
    }

}
