# ==========================================================================
# 
#       sound_ipaq.cdl
# 
#       eCos configuration data for the iPAQ audio device driver
# 
# ==========================================================================
# ####COPYRIGHTBEGIN####
#                                                                           
#  -------------------------------------------                              
#  The contents of this file are subject to the Red Hat eCos Public License 
#  Version 1.1 (the "License"); you may not use this file except in         
#  compliance with the License.  You may obtain a copy of the License at    
#  http://www.redhat.com/                                                   
#                                                                           
#  Software distributed under the License is distributed on an "AS IS"      
#  basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
#  License for the specific language governing rights and limitations under 
#  the License.                                                             
#                                                                           
#  The Original Code is eCos - Embedded Configurable Operating System,      
#  released September 30, 1998.                                             
#                                                                           
#  The Initial Developer of the Original Code is 3G Lab Ltd.
#  Portions created by 3G Lab are                                          
#  Copyright (C) 2001 3G Lab Ltd.
#  All Rights Reserved.                                                     
#  -------------------------------------------                              
#                                                                           
# ####COPYRIGHTEND####
# ==========================================================================
# #####DESCRIPTIONBEGIN####
# 
#  Author(s):    dominic.ostrowski@3glab.com
#  Contributors: dominic.ostrowski@3glab.com
#  Date:         2000-04-11
#  Purpose:      
#  Description:  Sound driver for the Compaq iPAQ
#               
# 
# ####DESCRIPTIONEND####
# 
# ==========================================================================


cdl_package CYGPKG_DEVS_SOUND_ARM_IPAQ {
	display		"Sound driver for iPAQ"
	include_dir	cyg/io
	requires	CYGPKG_IO
	requires	CYGFUN_KERNEL_API_C
	requires	CYGPKG_HAL_ARM_SA11X0_IPAQ
	description	"Sound driver for the iPAQ"
	compile		-library=libextras.a sound_ipaq.c

	cdl_component	CYGPKG_DEVS_SOUND_ARM_IPAQ_OPTIONS {
		display	"options"
		flavor	none
		no_define

		cdl_option	CYGDAT_DEVS_SOUND_ARM_IPAQ_NAME {
		    display	"Device name for the sound driver"
		    flavor	data
		    default_value	{"\"/dev/sound\""}
		    description	" This option specifies the name of the sound device"
		}

		cdl_option	CYGPKG_DEVS_SOUND_ARM_IPAQ_TESTS {
		    display	"Sound tests"
		    flavor	data
		    no_define
		    calculated	{ "tests/sound_test" }
		    description	"This option names the tests available for the sound driver"
		}
	}
}




